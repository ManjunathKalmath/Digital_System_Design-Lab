module mux_4x1();
input 
endmodule
